/*Copyright 2019-2021 T-Head Semiconductor Co., Ltd.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/

// &ModuleBeg; @25
module ct_idu_ir_vrt(
  dp_vrt_inst0_dst_vreg,
  dp_vrt_inst0_dstv_reg,
  dp_vrt_inst0_dstv_vld,
  dp_vrt_inst0_srcv0_reg,
  dp_vrt_inst0_srcv0_vld,
  dp_vrt_inst0_srcv1_reg,
  dp_vrt_inst0_srcv1_vld,
  dp_vrt_inst0_srcv2_vld,
  dp_vrt_inst0_srcvm_vld,
  dp_vrt_inst0_vmla,
  dp_vrt_inst1_dst_vreg,
  dp_vrt_inst1_dstv_reg,
  dp_vrt_inst1_dstv_vld,
  dp_vrt_inst1_srcv0_reg,
  dp_vrt_inst1_srcv0_vld,
  dp_vrt_inst1_srcv1_reg,
  dp_vrt_inst1_srcv1_vld,
  dp_vrt_inst1_srcv2_vld,
  dp_vrt_inst1_srcvm_vld,
  dp_vrt_inst1_vmla,
  dp_vrt_inst2_dst_vreg,
  dp_vrt_inst2_dstv_reg,
  dp_vrt_inst2_dstv_vld,
  dp_vrt_inst2_srcv0_reg,
  dp_vrt_inst2_srcv0_vld,
  dp_vrt_inst2_srcv1_reg,
  dp_vrt_inst2_srcv1_vld,
  dp_vrt_inst2_srcv2_vld,
  dp_vrt_inst2_srcvm_vld,
  dp_vrt_inst2_vmla,
  dp_vrt_inst3_dst_vreg,
  dp_vrt_inst3_dstv_reg,
  dp_vrt_inst3_dstv_vld,
  dp_vrt_inst3_srcv0_reg,
  dp_vrt_inst3_srcv0_vld,
  dp_vrt_inst3_srcv1_reg,
  dp_vrt_inst3_srcv1_vld,
  dp_vrt_inst3_srcv2_vld,
  dp_vrt_inst3_srcvm_vld,
  dp_vrt_inst3_vmla,
  rtu_idu_rt_recover_vreg,
  vrt_dp_inst01_srcv2_match,
  vrt_dp_inst02_srcv2_match,
  vrt_dp_inst03_srcv2_match,
  vrt_dp_inst0_rel_vreg,
  vrt_dp_inst0_srcv0_data,
  vrt_dp_inst0_srcv1_data,
  vrt_dp_inst0_srcv2_data,
  vrt_dp_inst0_srcvm_data,
  vrt_dp_inst12_srcv2_match,
  vrt_dp_inst13_srcv2_match,
  vrt_dp_inst1_rel_vreg,
  vrt_dp_inst1_srcv0_data,
  vrt_dp_inst1_srcv1_data,
  vrt_dp_inst1_srcv2_data,
  vrt_dp_inst1_srcvm_data,
  vrt_dp_inst23_srcv2_match,
  vrt_dp_inst2_rel_vreg,
  vrt_dp_inst2_srcv0_data,
  vrt_dp_inst2_srcv1_data,
  vrt_dp_inst2_srcv2_data,
  vrt_dp_inst2_srcvm_data,
  vrt_dp_inst3_rel_vreg,
  vrt_dp_inst3_srcv0_data,
  vrt_dp_inst3_srcv1_data,
  vrt_dp_inst3_srcv2_data,
  vrt_dp_inst3_srcvm_data
);

// &Ports; @26
input   [5  :0]  dp_vrt_inst0_dst_vreg;    
input   [5  :0]  dp_vrt_inst0_dstv_reg;    
input            dp_vrt_inst0_dstv_vld;    
input   [5  :0]  dp_vrt_inst0_srcv0_reg;   
input            dp_vrt_inst0_srcv0_vld;   
input   [5  :0]  dp_vrt_inst0_srcv1_reg;   
input            dp_vrt_inst0_srcv1_vld;   
input            dp_vrt_inst0_srcv2_vld;   
input            dp_vrt_inst0_srcvm_vld;   
input            dp_vrt_inst0_vmla;        
input   [5  :0]  dp_vrt_inst1_dst_vreg;    
input   [5  :0]  dp_vrt_inst1_dstv_reg;    
input            dp_vrt_inst1_dstv_vld;    
input   [5  :0]  dp_vrt_inst1_srcv0_reg;   
input            dp_vrt_inst1_srcv0_vld;   
input   [5  :0]  dp_vrt_inst1_srcv1_reg;   
input            dp_vrt_inst1_srcv1_vld;   
input            dp_vrt_inst1_srcv2_vld;   
input            dp_vrt_inst1_srcvm_vld;   
input            dp_vrt_inst1_vmla;        
input   [5  :0]  dp_vrt_inst2_dst_vreg;    
input   [5  :0]  dp_vrt_inst2_dstv_reg;    
input            dp_vrt_inst2_dstv_vld;    
input   [5  :0]  dp_vrt_inst2_srcv0_reg;   
input            dp_vrt_inst2_srcv0_vld;   
input   [5  :0]  dp_vrt_inst2_srcv1_reg;   
input            dp_vrt_inst2_srcv1_vld;   
input            dp_vrt_inst2_srcv2_vld;   
input            dp_vrt_inst2_srcvm_vld;   
input            dp_vrt_inst2_vmla;        
input   [5  :0]  dp_vrt_inst3_dst_vreg;    
input   [5  :0]  dp_vrt_inst3_dstv_reg;    
input            dp_vrt_inst3_dstv_vld;    
input   [5  :0]  dp_vrt_inst3_srcv0_reg;   
input            dp_vrt_inst3_srcv0_vld;   
input   [5  :0]  dp_vrt_inst3_srcv1_reg;   
input            dp_vrt_inst3_srcv1_vld;   
input            dp_vrt_inst3_srcv2_vld;   
input            dp_vrt_inst3_srcvm_vld;   
input            dp_vrt_inst3_vmla;        
input   [191:0]  rtu_idu_rt_recover_vreg;  
output           vrt_dp_inst01_srcv2_match; 
output           vrt_dp_inst02_srcv2_match; 
output           vrt_dp_inst03_srcv2_match; 
output  [6  :0]  vrt_dp_inst0_rel_vreg;    
output  [8  :0]  vrt_dp_inst0_srcv0_data;  
output  [8  :0]  vrt_dp_inst0_srcv1_data;  
output  [9  :0]  vrt_dp_inst0_srcv2_data;  
output  [8  :0]  vrt_dp_inst0_srcvm_data;  
output           vrt_dp_inst12_srcv2_match; 
output           vrt_dp_inst13_srcv2_match; 
output  [6  :0]  vrt_dp_inst1_rel_vreg;    
output  [8  :0]  vrt_dp_inst1_srcv0_data;  
output  [8  :0]  vrt_dp_inst1_srcv1_data;  
output  [9  :0]  vrt_dp_inst1_srcv2_data;  
output  [8  :0]  vrt_dp_inst1_srcvm_data;  
output           vrt_dp_inst23_srcv2_match; 
output  [6  :0]  vrt_dp_inst2_rel_vreg;    
output  [8  :0]  vrt_dp_inst2_srcv0_data;  
output  [8  :0]  vrt_dp_inst2_srcv1_data;  
output  [9  :0]  vrt_dp_inst2_srcv2_data;  
output  [8  :0]  vrt_dp_inst2_srcvm_data;  
output  [6  :0]  vrt_dp_inst3_rel_vreg;    
output  [8  :0]  vrt_dp_inst3_srcv0_data;  
output  [8  :0]  vrt_dp_inst3_srcv1_data;  
output  [9  :0]  vrt_dp_inst3_srcv2_data;  
output  [8  :0]  vrt_dp_inst3_srcvm_data;  

// &Regs; @27

// &Wires; @28
wire             vrt_dp_inst01_srcv2_match; 
wire             vrt_dp_inst02_srcv2_match; 
wire             vrt_dp_inst03_srcv2_match; 
wire    [6  :0]  vrt_dp_inst0_rel_vreg;    
wire    [8  :0]  vrt_dp_inst0_srcv0_data;  
wire    [8  :0]  vrt_dp_inst0_srcv1_data;  
wire    [9  :0]  vrt_dp_inst0_srcv2_data;  
wire    [8  :0]  vrt_dp_inst0_srcvm_data;  
wire             vrt_dp_inst12_srcv2_match; 
wire             vrt_dp_inst13_srcv2_match; 
wire    [6  :0]  vrt_dp_inst1_rel_vreg;    
wire    [8  :0]  vrt_dp_inst1_srcv0_data;  
wire    [8  :0]  vrt_dp_inst1_srcv1_data;  
wire    [9  :0]  vrt_dp_inst1_srcv2_data;  
wire    [8  :0]  vrt_dp_inst1_srcvm_data;  
wire             vrt_dp_inst23_srcv2_match; 
wire    [6  :0]  vrt_dp_inst2_rel_vreg;    
wire    [8  :0]  vrt_dp_inst2_srcv0_data;  
wire    [8  :0]  vrt_dp_inst2_srcv1_data;  
wire    [9  :0]  vrt_dp_inst2_srcv2_data;  
wire    [8  :0]  vrt_dp_inst2_srcvm_data;  
wire    [6  :0]  vrt_dp_inst3_rel_vreg;    
wire    [8  :0]  vrt_dp_inst3_srcv0_data;  
wire    [8  :0]  vrt_dp_inst3_srcv1_data;  
wire    [9  :0]  vrt_dp_inst3_srcv2_data;  
wire    [8  :0]  vrt_dp_inst3_srcvm_data;  


// &Force("bus","dp_rt_dep_info",DEP_WIDTH-1,0); @57
// &Instance("gated_clk_cell", "x_vrt_gated_clk"); @73
// &Connect(.clk_in      (forever_cpuclk), @74
//          .external_en (1'b0), @75
//          .global_en   (cp0_yy_clk_en), @76
//          .module_en   (cp0_idu_icg_en), @77
//          .local_en    (vrt_clk_en), @78
//          .clk_out     (vrt_top_clk)); @79
// &ConnRule(s/^x_/reg_0_/); @85
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_0"); @86
// &Connect(.forever_cpuclk(vrt_top_clk)); @87
// &ConnRule(s/^x_/reg_1_/); @88
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_1"); @89
// &Connect(.forever_cpuclk(vrt_top_clk)); @90
// &ConnRule(s/^x_/reg_2_/); @91
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_2"); @92
// &Connect(.forever_cpuclk(vrt_top_clk)); @93
// &ConnRule(s/^x_/reg_3_/); @94
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_3"); @95
// &Connect(.forever_cpuclk(vrt_top_clk)); @96
// &ConnRule(s/^x_/reg_4_/); @97
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_4"); @98
// &Connect(.forever_cpuclk(vrt_top_clk)); @99
// &ConnRule(s/^x_/reg_5_/); @100
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_5"); @101
// &Connect(.forever_cpuclk(vrt_top_clk)); @102
// &ConnRule(s/^x_/reg_6_/); @103
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_6"); @104
// &Connect(.forever_cpuclk(vrt_top_clk)); @105
// &ConnRule(s/^x_/reg_7_/); @106
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_7"); @107
// &Connect(.forever_cpuclk(vrt_top_clk)); @108
// &ConnRule(s/^x_/reg_8_/); @109
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_8"); @110
// &Connect(.forever_cpuclk(vrt_top_clk)); @111
// &ConnRule(s/^x_/reg_9_/); @112
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_9"); @113
// &Connect(.forever_cpuclk(vrt_top_clk)); @114
// &ConnRule(s/^x_/reg_10_/); @115
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_10"); @116
// &Connect(.forever_cpuclk(vrt_top_clk)); @117
// &ConnRule(s/^x_/reg_11_/); @118
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_11"); @119
// &Connect(.forever_cpuclk(vrt_top_clk)); @120
// &ConnRule(s/^x_/reg_12_/); @121
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_12"); @122
// &Connect(.forever_cpuclk(vrt_top_clk)); @123
// &ConnRule(s/^x_/reg_13_/); @124
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_13"); @125
// &Connect(.forever_cpuclk(vrt_top_clk)); @126
// &ConnRule(s/^x_/reg_14_/); @127
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_14"); @128
// &Connect(.forever_cpuclk(vrt_top_clk)); @129
// &ConnRule(s/^x_/reg_15_/); @130
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_15"); @131
// &Connect(.forever_cpuclk(vrt_top_clk)); @132
// &ConnRule(s/^x_/reg_16_/); @133
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_16"); @134
// &Connect(.forever_cpuclk(vrt_top_clk)); @135
// &ConnRule(s/^x_/reg_17_/); @136
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_17"); @137
// &Connect(.forever_cpuclk(vrt_top_clk)); @138
// &ConnRule(s/^x_/reg_18_/); @139
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_18"); @140
// &Connect(.forever_cpuclk(vrt_top_clk)); @141
// &ConnRule(s/^x_/reg_19_/); @142
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_19"); @143
// &Connect(.forever_cpuclk(vrt_top_clk)); @144
// &ConnRule(s/^x_/reg_20_/); @145
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_20"); @146
// &Connect(.forever_cpuclk(vrt_top_clk)); @147
// &ConnRule(s/^x_/reg_21_/); @148
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_21"); @149
// &Connect(.forever_cpuclk(vrt_top_clk)); @150
// &ConnRule(s/^x_/reg_22_/); @151
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_22"); @152
// &Connect(.forever_cpuclk(vrt_top_clk)); @153
// &ConnRule(s/^x_/reg_23_/); @154
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_23"); @155
// &Connect(.forever_cpuclk(vrt_top_clk)); @156
// &ConnRule(s/^x_/reg_24_/); @157
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_24"); @158
// &Connect(.forever_cpuclk(vrt_top_clk)); @159
// &ConnRule(s/^x_/reg_25_/); @160
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_25"); @161
// &Connect(.forever_cpuclk(vrt_top_clk)); @162
// &ConnRule(s/^x_/reg_26_/); @163
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_26"); @164
// &Connect(.forever_cpuclk(vrt_top_clk)); @165
// &ConnRule(s/^x_/reg_27_/); @166
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_27"); @167
// &Connect(.forever_cpuclk(vrt_top_clk)); @168
// &ConnRule(s/^x_/reg_28_/); @169
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_28"); @170
// &Connect(.forever_cpuclk(vrt_top_clk)); @171
// &ConnRule(s/^x_/reg_29_/); @172
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_29"); @173
// &Connect(.forever_cpuclk(vrt_top_clk)); @174
// &ConnRule(s/^x_/reg_30_/); @175
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_30"); @176
// &Connect(.forever_cpuclk(vrt_top_clk)); @177
// &ConnRule(s/^x_/reg_31_/); @178
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_31"); @179
// &Connect(.forever_cpuclk(vrt_top_clk)); @180
// &ConnRule(s/^x_/reg_32_/); @181
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_32"); @182
// &Connect(.forever_cpuclk(vrt_top_clk)); @183
// &ConnRule(s/^x_/reg_33_/); @184
// &Instance("ct_idu_dep_vreg_srcv2_entry","x_ct_idu_ir_vrt_entry_vreg_33"); @185
// &Connect(.forever_cpuclk(vrt_top_clk)); @186
// &ConnRule(s/^x_num/dp_vrt_inst0_dstv_reg_lsb/); @314
// &Instance("ct_rtu_expand_32","x_ct_rtu_expand_32_dp_vrt_inst0_dstv_reg_lsb"); @315
// &ConnRule(s/^x_num/dp_vrt_inst1_dstv_reg_lsb/); @316
// &Instance("ct_rtu_expand_32","x_ct_rtu_expand_32_dp_vrt_inst1_dstv_reg_lsb"); @317
// &ConnRule(s/^x_num/dp_vrt_inst2_dstv_reg_lsb/); @318
// &Instance("ct_rtu_expand_32","x_ct_rtu_expand_32_dp_vrt_inst2_dstv_reg_lsb"); @319
// &ConnRule(s/^x_num/dp_vrt_inst3_dstv_reg_lsb/); @320
// &Instance("ct_rtu_expand_32","x_ct_rtu_expand_32_dp_vrt_inst3_dstv_reg_lsb"); @321
// &CombBeg; @537
// &CombEnd; @548
// &CombBeg; @549
// &CombEnd; @560
// &CombBeg; @561
// &CombEnd; @572
// &CombBeg; @573
// &CombEnd; @584
// &CombBeg; @585
// &CombEnd; @596
// &CombBeg; @597
// &CombEnd; @608
// &CombBeg; @609
// &CombEnd; @620
// &CombBeg; @621
// &CombEnd; @632
// &CombBeg; @633
// &CombEnd; @644
// &CombBeg; @645
// &CombEnd; @656
// &CombBeg; @657
// &CombEnd; @668
// &CombBeg; @669
// &CombEnd; @680
// &CombBeg; @681
// &CombEnd; @692
// &CombBeg; @693
// &CombEnd; @704
// &CombBeg; @705
// &CombEnd; @716
// &CombBeg; @717
// &CombEnd; @728
// &CombBeg; @729
// &CombEnd; @740
// &CombBeg; @741
// &CombEnd; @752
// &CombBeg; @753
// &CombEnd; @764
// &CombBeg; @765
// &CombEnd; @776
// &CombBeg; @777
// &CombEnd; @788
// &CombBeg; @789
// &CombEnd; @800
// &CombBeg; @801
// &CombEnd; @812
// &CombBeg; @813
// &CombEnd; @824
// &CombBeg; @825
// &CombEnd; @836
// &CombBeg; @837
// &CombEnd; @848
// &CombBeg; @849
// &CombEnd; @860
// &CombBeg; @861
// &CombEnd; @872
// &CombBeg; @873
// &CombEnd; @884
// &CombBeg; @885
// &CombEnd; @896
// &CombBeg; @897
// &CombEnd; @908
// &CombBeg; @909
// &CombEnd; @920
// &CombBeg; @921
// &CombEnd; @932
// &CombBeg; @933
// &CombEnd; @944
// &CombBeg; @988
// &CombEnd; @1026
// &CombBeg; @1039
// &CombEnd; @1077
// &CombBeg; @1090
// &CombEnd; @1128
// &CombBeg; @1167
// &CombEnd; @1205
// &CombBeg; @1222
// &CombEnd; @1235
// &CombBeg; @1238
// &CombEnd; @1276
// &CombBeg; @1295
// &CombEnd; @1308
// &CombBeg; @1311
// &CombEnd; @1349
// &CombBeg; @1368
// &CombEnd; @1389
// &CombBeg; @1408
// &CombEnd; @1421
// &CombBeg; @1439
// &CombEnd; @1446
// &CombBeg; @1452
// &CombEnd; @1490
// &CombBeg; @1512
// &CombEnd; @1530
// &CombBeg; @1533
// &CombEnd; @1571
// &CombBeg; @1592
// &CombEnd; @1610
// &CombBeg; @1613
// &CombEnd; @1651
// &CombBeg; @1672
// &CombEnd; @1704
// &CombBeg; @1725
// &CombEnd; @1743
// &CombBeg; @1760
// &CombEnd; @1769
// &CombBeg; @1775
// &CombEnd; @1813
// &CombBeg; @1842
// &CombEnd; @1865
// &CombBeg; @1868
// &CombEnd; @1906
// &CombBeg; @1932
// &CombEnd; @1955
// &CombBeg; @1958
// &CombEnd; @1996
// &CombBeg; @2022
// &CombEnd; @2067
// &CombBeg; @2093
// &CombEnd; @2116
// &CombBeg; @2137
// &CombEnd; @2148
// &Force("input","dp_vrt_inst0_dst_vreg"); @2151
// &Force("input","dp_vrt_inst0_dstv_reg"); @2152
// &Force("input","dp_vrt_inst0_dstv_vld"); @2153
// &Force("input","dp_vrt_inst0_srcv0_reg"); @2154
// &Force("input","dp_vrt_inst0_srcv0_vld"); @2155
// &Force("input","dp_vrt_inst0_srcv1_reg"); @2156
// &Force("input","dp_vrt_inst0_srcv1_vld"); @2157
// &Force("input","dp_vrt_inst0_srcv2_vld"); @2158
// &Force("input","dp_vrt_inst0_srcvm_vld"); @2159
// &Force("input","dp_vrt_inst0_vmla"); @2160
// &Force("input","dp_vrt_inst1_dst_vreg"); @2161
// &Force("input","dp_vrt_inst1_dstv_reg"); @2162
// &Force("input","dp_vrt_inst1_dstv_vld"); @2163
// &Force("input","dp_vrt_inst1_srcv0_reg"); @2164
// &Force("input","dp_vrt_inst1_srcv0_vld"); @2165
// &Force("input","dp_vrt_inst1_srcv1_reg"); @2166
// &Force("input","dp_vrt_inst1_srcv1_vld"); @2167
// &Force("input","dp_vrt_inst1_srcv2_vld"); @2168
// &Force("input","dp_vrt_inst1_srcvm_vld"); @2169
// &Force("input","dp_vrt_inst1_vmla"); @2170
// &Force("input","dp_vrt_inst2_dst_vreg"); @2171
// &Force("input","dp_vrt_inst2_dstv_reg"); @2172
// &Force("input","dp_vrt_inst2_dstv_vld"); @2173
// &Force("input","dp_vrt_inst2_srcv0_reg"); @2174
// &Force("input","dp_vrt_inst2_srcv0_vld"); @2175
// &Force("input","dp_vrt_inst2_srcv1_reg"); @2176
// &Force("input","dp_vrt_inst2_srcv1_vld"); @2177
// &Force("input","dp_vrt_inst2_srcv2_vld"); @2178
// &Force("input","dp_vrt_inst2_srcvm_vld"); @2179
// &Force("input","dp_vrt_inst2_vmla"); @2180
// &Force("input","dp_vrt_inst3_dst_vreg"); @2181
// &Force("input","dp_vrt_inst3_dstv_reg"); @2182
// &Force("input","dp_vrt_inst3_dstv_vld"); @2183
// &Force("input","dp_vrt_inst3_srcv0_reg"); @2184
// &Force("input","dp_vrt_inst3_srcv0_vld"); @2185
// &Force("input","dp_vrt_inst3_srcv1_reg"); @2186
// &Force("input","dp_vrt_inst3_srcv1_vld"); @2187
// &Force("input","dp_vrt_inst3_srcv2_vld"); @2188
// &Force("input","dp_vrt_inst3_srcvm_vld"); @2189
// &Force("input","dp_vrt_inst3_vmla"); @2190
// &Force("input","rtu_idu_rt_recover_vreg"); @2191

// &Force("bus","dp_vrt_inst0_dst_vreg",5,0); @2193
// &Force("bus","dp_vrt_inst0_dstv_reg",5,0); @2194
// &Force("bus","dp_vrt_inst0_srcv0_reg",5,0); @2195
// &Force("bus","dp_vrt_inst0_srcv1_reg",5,0); @2196
// &Force("bus","dp_vrt_inst1_dst_vreg",5,0); @2197
// &Force("bus","dp_vrt_inst1_dstv_reg",5,0); @2198
// &Force("bus","dp_vrt_inst1_srcv0_reg",5,0); @2199
// &Force("bus","dp_vrt_inst1_srcv1_reg",5,0); @2200
// &Force("bus","dp_vrt_inst2_dst_vreg",5,0); @2201
// &Force("bus","dp_vrt_inst2_dstv_reg",5,0); @2202
// &Force("bus","dp_vrt_inst2_srcv0_reg",5,0); @2203
// &Force("bus","dp_vrt_inst2_srcv1_reg",5,0); @2204
// &Force("bus","dp_vrt_inst3_dst_vreg",5,0); @2205
// &Force("bus","dp_vrt_inst3_dstv_reg",5,0); @2206
// &Force("bus","dp_vrt_inst3_srcv0_reg",5,0); @2207
// &Force("bus","dp_vrt_inst3_srcv1_reg",5,0); @2208
// &Force("bus","rtu_idu_rt_recover_vreg",191,0); @2209

assign vrt_dp_inst01_srcv2_match    = 1'b0;
assign vrt_dp_inst02_srcv2_match    = 1'b0;
assign vrt_dp_inst03_srcv2_match    = 1'b0;
assign vrt_dp_inst0_rel_vreg[6:0]   = 7'b0;
assign vrt_dp_inst0_srcv0_data[8:0] = 9'b100000011;
assign vrt_dp_inst0_srcv1_data[8:0] = 9'b100000011;
assign vrt_dp_inst0_srcv2_data[9:0] = 10'b1000000111;
assign vrt_dp_inst0_srcvm_data[8:0] = 9'b100000011;
assign vrt_dp_inst12_srcv2_match    = 1'b0;
assign vrt_dp_inst13_srcv2_match    = 1'b0;
assign vrt_dp_inst1_rel_vreg[6:0]   = 7'b0;
assign vrt_dp_inst1_srcv0_data[8:0] = 9'b100000011;
assign vrt_dp_inst1_srcv1_data[8:0] = 9'b100000011;
assign vrt_dp_inst1_srcv2_data[9:0] = 10'b1000000111;
assign vrt_dp_inst1_srcvm_data[8:0] = 9'b100000011;
assign vrt_dp_inst23_srcv2_match    = 1'b0;
assign vrt_dp_inst2_rel_vreg[6:0]   = 7'b0;
assign vrt_dp_inst2_srcv0_data[8:0] = 9'b100000011;
assign vrt_dp_inst2_srcv1_data[8:0] = 9'b100000011;
assign vrt_dp_inst2_srcv2_data[9:0] = 10'b1000000111;
assign vrt_dp_inst2_srcvm_data[8:0] = 9'b100000011;
assign vrt_dp_inst3_rel_vreg[6:0]   = 7'b0;
assign vrt_dp_inst3_srcv0_data[8:0] = 9'b100000011;
assign vrt_dp_inst3_srcv1_data[8:0] = 9'b100000011;
assign vrt_dp_inst3_srcv2_data[9:0] = 10'b1000000111;
assign vrt_dp_inst3_srcvm_data[8:0] = 9'b100000011;


// &ModuleEnd; @2240
endmodule


